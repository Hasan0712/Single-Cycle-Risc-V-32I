module register_tb ();
    reg [31:0]data_tb;
    reg clk;
    reg reset;
    reg enable;
    reg [4:0]rs1addr;
    reg [4:0]rs2addr;
    reg [4:0]rdaddr;
    wire [31:0] opa;
    wire [31:0] opb;
    









endmodule